library vunit_lib;
context vunit_lib.vunit_context;
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;


entity tb_top is
  generic (runner_cfg : string);
end entity;

architecture tb of tb_top is

  signal LED_G : std_logic;
  signal LED_R : std_logic;

  signal cpld_clk : std_logic;
    
    -----------------------------------------------------------------
    -- M65 Serial monitor interface
    -----------------------------------------------------------------    
    -- UART pins on the JB1 JTAG connector
  signal te_uart_tx : std_logic;
  signal te_uart_rx : std_logic;

    -- The UART pins on the Xilinx FPGA
  signal dbg_uart_tx : std_logic;
  signal dbg_uart_rx : std_logic;

    -----------------------------------------------------------------
    -- MAX10 own debug UART interface
    -----------------------------------------------------------------
    -- (overloads external uSD card interface, so we have to tri-state
    --  it).
  signal m_tx : std_logic := 'Z';
  signal m_rx : std_logic;
    
    -----------------------------------------------------------------
    -- Motherboard dip-switches: All off by default
    -----------------------------------------------------------------
  signal cpld_cfg0 : std_logic := '0';
  signal cpld_cfg1 : std_logic := '0';
  signal cpld_cfg2 : std_logic := '0';
  signal cpld_cfg3 : std_logic := '0';

    -----------------------------------------------------------------
    -- J21 GPIO interface
    -----------------------------------------------------------------
  signal J21 : std_logic_vector(11 downto 0) := (others => '0');
    
    -----------------------------------------------------------------
   -- Xilinx FPGA JTAG interface
    -----------------------------------------------------------------
    -- FPGA pins
  signal fpga_tck : std_logic;
  signal fpga_tdo : std_logic;
  signal fpga_tdi : std_logic;
  signal fpga_tms : std_logic;
    -- TE0790 pins
  signal te_tck : std_logic;
  signal te_tdo : std_logic;
  signal te_tdi : std_logic;
  signal te_tms : std_logic;
        
    -----------------------------------------------------------------
    -- Xilinx FPGA configuration control
    -----------------------------------------------------------------
  signal fpga_prog_b : std_logic := 'Z';
  signal fpga_init : std_logic := 'Z';
  signal fpga_done : std_logic;   
    
    -----------------------------------------------------------------
    -- Xilinx FPGA communications channel
    -----------------------------------------------------------------
  signal xilinx_sync : std_logic;
  signal xilinx_tx : std_logic;
  signal xilinx_rx : std_logic := '1';
    
    -----------------------------------------------------------------
    -- 5V Power rail control
    -----------------------------------------------------------------
  signal en_5v_joy_n : std_logic := '0';

    -----------------------------------------------------------------
    -- Keyboard connector
    -----------------------------------------------------------------
    -- pins connecting to xilinx fpga
  signal kb_tdo : std_logic;
  signal kb_tdi : std_logic;
  signal kb_tck : std_logic;
  signal kb_tms : std_logic;
  signal kb_jtagen : std_logic;
  signal kb_io1 : std_logic;
  signal kb_io2 : std_logic;
  signal kb_io3 : std_logic;
    -- pins connecting to actual keyboard
  signal k_tdo : std_logic;
  signal k_tdi : std_logic;
  signal k_tck : std_logic;
  signal k_tms : std_logic;
  signal k_jtagen : std_logic;
  signal k_io1 : std_logic;
  signal k_io2 : std_logic;
  signal k_io3 : std_logic;

    -----------------------------------------------------------------
    -- Reset button
    -----------------------------------------------------------------
  signal reset_btn : std_logic;
  signal blue_wire : std_logic;

  signal SCAN_OUT    : std_logic_vector(9 downto 0);
  signal SCAN_IN    : std_logic_vector(7 downto 0);
  
    -- A selection of keys to model
  signal key_f    : std_logic := '1'; -- Column 2, row 5
  signal key_o    : std_logic := '1'; -- Column 4, row 6,
  signal key_RETURN    : std_logic := '1'; -- Column 0, row 1
  signal key_UP    : std_logic := '1'; -- Colum 0, row 7 + Column 6, row 4 (RSHIFT)
  signal key_DOWN    : std_logic := '1'; -- Column 0, row 7

  signal mk1_KIO8    : std_logic;
  signal mk1_KIO9    : std_logic;
  signal mk1_KIO10    : std_logic;

  signal mk2_KIO8    : std_logic;
  signal mk2_KIO9    : std_logic;
  signal mk2_KIO10    : std_logic;
  
  signal KIO8    : std_logic;
  signal KIO9    : std_logic;
  signal KIO10    : std_logic;
    
  signal KEY_RESTORE    : std_logic;
  
  signal LED_R0    : std_logic;
  signal LED_G0    : std_logic;
  signal LED_B0    : std_logic;
  
  signal LED_R1    : std_logic;
  signal LED_G1    : std_logic;
  signal LED_B1    : std_logic;
  
  signal LED_R2    : std_logic;
  signal LED_G2    : std_logic;
  signal LED_B2    : std_logic;
  
  signal LED_R3    : std_logic;
  signal LED_G3    : std_logic;
  signal LED_B3    : std_logic;
  
  signal LED_SHIFT    : std_logic;
  signal LED_CAPS    : std_logic;
      
    -----------------------------------------------------------------
    -- VGA VDAC low-power switch
    -----------------------------------------------------------------
  signal vdac_psave_n : std_logic := '1';

  -- High if we are simulating a MK-I keyboard being connected,
  -- or low if simulating a MK-II keyboard being connected.
  signal mk1_connected : std_logic := '1';
  
begin

  -- Simulation can select which keyboard type is connected
  process (mk1_connected) is
  begin
    if mk1_connected = '1' then
      -- MK-I keyboard connected
      mk1_KIO8 <= kb_io1;
      mk1_KIO9 <= kb_io2;
      kb_io3 <= mk1_KIO10;
    else
      -- MK-II keyboard connected
      -- This is tricker, as we have to make two-way connection
      -- for SDA (KIO8) at least.
      -- XXX Not implemented
      kb_io3 <= '0';
    end if;
  end process;
    
  
  mk1_keyboard0: entity work.keyboard
    port map (
      SCAN_OUT => SCAN_OUT,
      SCAN_IN => SCAN_IN,

      -- A selection of keys to model
      key_f => key_f ,
      key_o => key_o ,
      key_RETURN => key_RETURN ,
      key_UP => key_UP ,
      key_DOWN => key_DOWN 
      
      );
  
  mk1_cpld0: entity work.keyboard_cpld
    port map (
      KIO8 => mk1_KIO8 ,
      KIO9 => mk1_KIO9 ,
      KIO10 => mk1_KIO10 ,
    
      SCAN_OUT	=> SCAN_OUT,
      SCAN_IN	=> SCAN_IN,
    
    
      KEY_RESTORE => KEY_RESTORE,
    
      LED_R0           	=> LED_R0,
      LED_G0           	=> LED_G0,
      LED_B0           	=> LED_B0,
   
      LED_R1           	=> LED_R1,
      LED_G1           	=> LED_G1,
      LED_B1           	=> LED_B1,
    
      LED_R2           	=> LED_R2,
      LED_G2           	=> LED_G2,
      LED_B2           	=> LED_B2,
    
      LED_R3           	=> LED_R3,
      LED_G3           	=> LED_G3,
      LED_B3           	=> LED_B3,
    
      LED_SHIFT           => LED_SHIFT,
      LED_CAPS            => LED_CAPS
      );
  
  top0: entity work.top
    port map (

      LED_G => LED_G,
      LED_R => LED_R,

      cpld_clk => cpld_clk,
    
    -----------------------------------------------------------------
    -- M65 Serial monitor interface
    -----------------------------------------------------------------    
    -- UART pins on the JB1 JTAG connector
      te_uart_tx => te_uart_tx,
      te_uart_rx => te_uart_rx,

    -- The UART pins on the Xilinx FPGA
      dbg_uart_tx => dbg_uart_tx,
      dbg_uart_rx => dbg_uart_rx,

    -----------------------------------------------------------------
    -- MAX10 own debug UART interface
    -----------------------------------------------------------------
    -- (overloads external uSD card interface, so we have to tri-state
    --  it).
      m_tx => m_tx,
      m_rx => m_rx,
    
    -----------------------------------------------------------------
    -- Motherboard dip-switches
    -----------------------------------------------------------------
      cpld_cfg0 => cpld_cfg0,
      cpld_cfg1 => cpld_cfg1,
      cpld_cfg2 => cpld_cfg2,
      cpld_cfg3 => cpld_cfg3,

    -----------------------------------------------------------------
    -- J21 GPIO interface
    -----------------------------------------------------------------
      J21 => J21,
    
    -----------------------------------------------------------------
   -- Xilinx FPGA JTAG interface
    -----------------------------------------------------------------
    -- FPGA pins
      fpga_tck => fpga_tck,
      fpga_tdo => fpga_tdo,
      fpga_tdi => fpga_tdi,
      fpga_tms => fpga_tms,
    -- TE0790 pins
      te_tck => te_tck,
      te_tdo => te_tdo,
      te_tdi => te_tdi,
      te_tms => te_tms,
        
    -----------------------------------------------------------------
    -- Xilinx FPGA configuration control
    -----------------------------------------------------------------
      fpga_prog_b => fpga_prog_b,
      fpga_init => fpga_init,
      fpga_done => fpga_done,
    
    -----------------------------------------------------------------
    -- Xilinx FPGA communications channel
    -----------------------------------------------------------------
      xilinx_sync => xilinx_sync,
      xilinx_tx => xilinx_tx,
      xilinx_rx => xilinx_rx,
    
    -----------------------------------------------------------------
    -- 5V Power rail control
    -----------------------------------------------------------------
      en_5v_joy_n => en_5v_joy_n,

    -----------------------------------------------------------------
    -- Keyboard connector
    -----------------------------------------------------------------
    -- pins connecting to xilinx fpga
      kb_tdo => kb_tdo,
      kb_tdi => kb_tdi,
      kb_tck => kb_tck,
      kb_tms => kb_tms,
      kb_jtagen => kb_jtagen,
      kb_io1 => kb_io1,
      kb_io2 => kb_io2,
      kb_io3 => kb_io3,
    -- pins connecting to actual keyboard
      k_tdo => k_tdo,
      k_tdi => k_tdi,
      k_tck => k_tck,
      k_tms => k_tms,
      k_jtagen => k_jtagen,
      k_io1 => k_io1,
      k_io2 => k_io2,
      k_io3 => k_io3,

    -----------------------------------------------------------------
    -- Reset button
    -----------------------------------------------------------------
      reset_btn => reset_btn,
      blue_wire => blue_wire,

    -----------------------------------------------------------------
    -- VGA VDAC low-power switch
    -----------------------------------------------------------------
      vdac_psave_n => vdac_psave_n
    
      );
   
  main : process
  begin
    test_runner_setup(runner, runner_cfg);
        
    while test_suite loop

      if run("MAX10 relays MK-I keyboard traffic to main FPGA") then
        assert false report "not implemented";
      end if;
    end loop;
    test_runner_cleanup(runner);
  end process;
end architecture;
