
module intclock (
	oscena,
	clkout);	

	input		oscena;
	output		clkout;
endmodule
