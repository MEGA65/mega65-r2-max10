
module intclock (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
